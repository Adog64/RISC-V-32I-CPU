module CPU ();
    wire[4:0] Q0, Q1, Q2;
    wire[11:0] Q4;
    wire[31:0] Q5, Q6, Q7, Q8, Q9, Q10, Q11, Q12, Q13, Q14, Q15, Q16;
    
    
endmodule